library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cla_16bit is 
port ( a : in STD_LOGIC_VECTOR (15 downto 0);
b : 