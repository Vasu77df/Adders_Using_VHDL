LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY fourbit_cla_t IS
END fourbit_cla_t;
 
ARCHITECTURE behavior OF fourbit_cla_t IS
 
-- Component Declaration for the Unit Under Test (UUT)
 
COMPONENT cla
PORT(
a : IN std_logic_vector(3 downto 0);
b : IN std_logic_vector(3 downto 0);
cin : IN std_logic;
s : OUT std_logic_vector(3 downto 0);
cout : OUT std_logic
);
END COMPONENT;
 
--Inputs
signal a : std_logic_vector(3 downto 0) := (others => '0');
signal b : std_logic_vector(3 downto 0) := (others => '0');
signal cin : std_logic := '0';
 
--Outputs
signal s : std_logic_vector(3 downto 0);
signal cout : std_logic;
 
BEGIN
 
-- Instantiate the Unit Under Test (UUT)
uut: cla PORT MAP (
a => a,
b => b,
cin => cin,
s => s,
cout => cout
);
 
-- Stimulus process
stim_proc: process
begin
-- hold reset state for 100 ns.
wait for 10 ns;
 
a <= "1111";
b <= "1111";
cin <= '1';
 
wait for 10 ns;
a <= "1010";
b <= "0111";
cin <= '0';
 
wait for 10 ns;
 
a <= "1000";
b <= "1001";
cin <= '0';
 
wait;
 
end process;
 
END;
