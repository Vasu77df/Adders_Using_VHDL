library ieee;
use ieee.std_logic_1164.all;

entity rca_thirtytwo_t is
end rca_thirtytwo_t;

architecture behav of rca_thirtytwo_t is 

COMPONENT rca_thirtytwo
PORT(
a : IN std_logic_vector(31 downto 0);
b : IN std_logic_vector(31 downto 0);
cin : IN std_logic;
s : OUT std_logic_vector(31 downto 0);
cout : OUT std_logic
);
END COMPONENT;

--Inputs
signal a : std_logic_vector(31 downto 0) := (others => '0');
signal b : std_logic_vector(31 downto 0) := (others => '0');
signal cin : std_logic := '0';

--Outputs
signal s : std_logic_vector(31 downto 0);
signal cout : std_logic;

BEGIN 

uut: rca_thirtytwo PORT MAP (
a => a,
b => b,
cin => cin,
s => s,
cout => cout
);

stim_proc: process 
begin 

wait for 10 ns;
a <= "00000000000000000000011111111100"; -- A id number first four bits that is 2044 
b <= "00000000000000000001011101110011"; -- A id number first four bits that is 6003
cin <= '0';

wait for 10 ns;
a <= "00000000000001000010011110111100";
b <= "00000000000100001001011101110011";
cin <= '1';

wait for 10 ns;
a <= "00000000000001000100011111101100";
b <= "00000000001010000001010101110011";
cin <= '1';

wait;

end process;

END;